// Example code for an M0 AHBLite System
//  Iain McNally
//  ECS, University of Soutampton
//
// This module is an AHB-Lite Slave containing a RAM
//
// Number of addressable locations : 2**MEMWIDTH
// Size of each addressable location : 8 bits
// Supported transfer sizes : Word, Halfword, Byte
// Alignment of base address : Word aligned
//


module ahb_ram #(
  parameter MEMWIDTH = 8
)(
  //AHBLITE INTERFACE

    //Slave Select Signal
    input HSEL,
    //Global Signals
    input HCLK,
    input HRESETn,
    //Address, Control & Write Data
    input HREADY,
    input [31:0] HADDR,
    input [1:0] HTRANS,
    input HWRITE,
    input [2:0] HSIZE,
    input [31:0] HWDATA,
    // Transfer Response & Read Data
    output HREADYOUT,
    output [31:0] HRDATA

);

timeunit 1ns;
timeprecision 100ps;

  localparam No_Transfer = 2'b0;

// control signals are stored in registers
  logic write_enable, read_enable;
  logic [MEMWIDTH-2:0] word_address;
  logic [3:0] byte_select;

// Macro Cell Signals
  logic [31:0] HWDATA_RAM;
  wire  [31:0] HRDATA_RAM;
  
// Instantiation
  sram256x32 sram256x32_1 (
    .NRST(HRESETn),
    .CS(HCLK),
    .RD(read_enable),
    .WR(write_enable),
    .EN(1'b0),
    .AD({word_address, 2'b0}),
    .DI(HWDATA),
    .DO(HRDATA_RAM)
  );


// Generate the control signals in the address phase
  always_ff @(posedge HCLK, negedge HRESETn)
    if (! HRESETn )
      begin
        write_enable <= '0;
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
      end
    else if ( HREADY && HSEL && (HTRANS != No_Transfer) )
      begin
        write_enable <= HWRITE;
        read_enable <= ! HWRITE;
        word_address <= HADDR[MEMWIDTH:2];
        byte_select <= generate_byte_select( HSIZE, HADDR[1:0] );
     end
    else
      begin
        write_enable <= '0;
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
     end

//Act on control signals in the data phase

//Transfer Response
  assign HREADYOUT = '1; //Single cycle Write & Read. Zero Wait state operations

// decode byte select signals from the size and the lowest two address bits
  function logic [3:0] generate_byte_select( logic [2:0] size, logic [1:0] byte_adress );
    logic byte3, byte2, byte1, byte0;
    byte0 = size[1] || ( byte_adress == 0 );
    byte1 = size[1] || ( size[0] && ( byte_adress == 0 ) ) || ( byte_adress == 1 );
    byte2 = size[1] || ( byte_adress == 2 );
    byte3 = size[1] || ( size[0] && ( byte_adress == 2 ) ) || ( byte_adress == 3 );
    return { byte3, byte2, byte1, byte0 };
  endfunction

endmodule
