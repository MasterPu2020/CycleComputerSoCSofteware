assign resource_rom[ 0] = 104'hFFFFFFFFFFFFFFE07F03F81FC0; // File Name: template.png
