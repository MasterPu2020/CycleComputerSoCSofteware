assign location_rom[ 0] = 16'h0000;
assign location_rom[ 1] = 16'h0008;
assign location_rom[ 2] = 16'h0010;
assign location_rom[ 3] = 16'h0018;
assign location_rom[ 4] = 16'h0020;
assign location_rom[ 5] = 16'h0028;
assign location_rom[ 6] = 16'h0030;
assign location_rom[ 7] = 16'h0038;
assign location_rom[ 8] = 16'h0040;
assign location_rom[ 9] = 16'h0D00;
assign location_rom[10] = 16'h0D08;
assign location_rom[11] = 16'h0D10;
assign location_rom[12] = 16'h0D18;
assign location_rom[13] = 16'h0D20;
assign location_rom[14] = 16'h0D28;
assign location_rom[15] = 16'h0D30;
assign location_rom[16] = 16'h0D38;
assign location_rom[17] = 16'h0D40;
assign location_rom[18] = 16'h1A00;
assign location_rom[19] = 16'h1A08;
assign location_rom[20] = 16'h1A10;
assign location_rom[21] = 16'h1A18;
assign location_rom[22] = 16'h1A20;
assign location_rom[23] = 16'h1A28;
assign location_rom[24] = 16'h1A30;
assign location_rom[25] = 16'h1A38;
assign location_rom[26] = 16'h1A40;
assign location_rom[27] = 16'h2700;
assign location_rom[28] = 16'h3400;
assign location_rom[29] = 16'h3408;
assign location_rom[30] = 16'h3410;
assign location_rom[31] = 16'h3418;
