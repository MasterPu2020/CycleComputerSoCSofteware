assign resource_rom[ 0] = 104'h7EFFC3C3C3C3C3C3C3C3C3FF7E; // File Name: 0.png
assign resource_rom[ 1] = 104'hFF7E18181818181818181B1E1C; // File Name: 1.png
assign resource_rom[ 2] = 104'h7EFFFF0303037FFEC0C0C0FF7E; // File Name: 2.png
assign resource_rom[ 3] = 104'h7EFFFFC0C0C0FFFFC0C0C0FF7F; // File Name: 3.png
assign resource_rom[ 4] = 104'h40C0C0C0C0FEFFFFC3C3C3C3C3; // File Name: 4.png
assign resource_rom[ 5] = 104'h7EFFFFC0C0C0FFFF030303FF7F; // File Name: 5.png
assign resource_rom[ 6] = 104'h7EFFFFC3C3C3FFFF030303FF7F; // File Name: 6.png
assign resource_rom[ 7] = 104'h40C0C0C0C0C0C0C0C0C0C0FFFE; // File Name: 7.png
assign resource_rom[ 8] = 104'h7EFFC3C3C3C3FFFFC3C3C3FF7E; // File Name: 8.png
assign resource_rom[ 9] = 104'h7EFFFFC0C0C0FEFFC3C3C3FF7E; // File Name: 9.png
assign resource_rom[10] = 104'h3C665A5A663CE09C3C00000000; // File Name: candence1.png
assign resource_rom[11] = 104'h3C665A5A663C1C090F0E041F1F; // File Name: candence2.png
assign resource_rom[12] = 104'h00000018180000001818000000; // File Name: colon.png
assign resource_rom[13] = 104'h8282868606060C8C8C98181890; // File Name: distance1.png
assign resource_rom[14] = 104'h41416161606030313119181809; // File Name: distance2.png
assign resource_rom[15] = 104'h00181800000000000000000000; // File Name: dot.png
assign resource_rom[16] = 104'h00000000000000000000000000; // File Name: empty.png
assign resource_rom[17] = 104'h330B0F0B330303030200000000; // File Name: km1.png
assign resource_rom[18] = 104'h2B2B2B2B3F1F00000000000000; // File Name: km2.png
assign resource_rom[19] = 104'h330B0F0B330303030200000000; // File Name: kmh1.png
assign resource_rom[20] = 104'h2B2B2B2B3F1F00000000000000; // File Name: kmh2.png
assign resource_rom[21] = 104'h13131313131F03030300000000; // File Name: kmh3.png
assign resource_rom[22] = 104'h565656567E3E00000000000000; // File Name: mm1.png
assign resource_rom[23] = 104'h565656567E3E00000000000000; // File Name: mm2.png
assign resource_rom[24] = 104'h00000606060E1E360000000000; // File Name: rpm1.png
assign resource_rom[25] = 104'h0303838F9F93938F0000000000; // File Name: rpm2.png
assign resource_rom[26] = 104'h0000151515151F0F0000000000; // File Name: rpm3.png
assign resource_rom[27] = 104'h78C888183060407C183060C080; // File Name: speed1.png
assign resource_rom[28] = 104'h00000103060C183E060C18103F; // File Name: speed2.png
assign resource_rom[29] = 104'hE0F0180C06868686868C18F0E0; // File Name: timer1.png
assign resource_rom[30] = 104'h070F1830606767606030180F07; // File Name: timer2.png
assign resource_rom[31] = 104'hCCDCF8F8F8787070E0C0800000; // File Name: timeunit1.png
assign resource_rom[32] = 104'h73F7FFFFFF9E9EDFFFFFFF7F00; // File Name: timeunit2.png
assign resource_rom[33] = 104'h060E1F1F1F1F1F0F0703010000; // File Name: timeunit3.png
