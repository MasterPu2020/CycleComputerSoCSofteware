assign location_rom[ 0] = 16'h0000;
assign location_rom[ 1] = 16'h0800;
assign location_rom[ 2] = 16'h1000;
assign location_rom[ 3] = 16'h1800;
assign location_rom[ 4] = 16'h2000;
assign location_rom[ 5] = 16'h2800;
assign location_rom[ 6] = 16'h3000;
assign location_rom[ 7] = 16'h3800;
assign location_rom[ 8] = 16'h4000;
assign location_rom[ 9] = 16'h000D;
assign location_rom[10] = 16'h080D;
assign location_rom[11] = 16'h100D;
assign location_rom[12] = 16'h180D;
assign location_rom[13] = 16'h200D;
assign location_rom[14] = 16'h280D;
assign location_rom[15] = 16'h300D;
assign location_rom[16] = 16'h380D;
assign location_rom[17] = 16'h400D;
assign location_rom[18] = 16'h001A;
assign location_rom[19] = 16'h081A;
assign location_rom[20] = 16'h101A;
assign location_rom[21] = 16'h181A;
assign location_rom[22] = 16'h201A;
assign location_rom[23] = 16'h281A;
assign location_rom[24] = 16'h301A;
assign location_rom[25] = 16'h381A;
assign location_rom[26] = 16'h401A;
assign location_rom[27] = 16'h0027;
assign location_rom[28] = 16'h0034;
assign location_rom[29] = 16'h0834;
assign location_rom[30] = 16'h1034;
assign location_rom[31] = 16'h1834;
