assign location_rom[ 0] = 16'h1F0E;
assign location_rom[ 1] = 16'h1F16;
assign location_rom[ 2] = 16'h1F2A;
assign location_rom[ 3] = 16'h2C35;
assign location_rom[ 4] = 16'h1F35;
assign location_rom[ 5] = 16'h2C45;
assign location_rom[ 6] = 16'h1F45;
assign location_rom[ 7] = 16'h2C50;
assign location_rom[ 8] = 16'h1F50;
assign location_rom[ 9] = 16'h1F5E;
assign location_rom[10] = 16'h1F66;
assign location_rom[11] = 16'h1F6E;
assign location_rom[12] = 16'h1F3D;
assign location_rom[13] = 16'h3E0E;
assign location_rom[14] = 16'h3E16;
assign location_rom[15] = 16'h3E2A;
assign location_rom[16] = 16'h3E35;
assign location_rom[17] = 16'h3E45;
assign location_rom[18] = 16'h3E50;
assign location_rom[19] = 16'h3E3D;
