assign resource_rom[ 0] = 104'hE7E7E7E7E7E7E7E70000E7E7E7; // File Name: template.png
